package types;
  typedef logic [15:0] f16;  // 16 bit float point
  typedef logic [15:0] fx13;  // 13 bit fixed point
  typedef logic signed [15:0] i13;  // 13 bit integer
  typedef f16 vec3_f16[3];
  typedef f16 vec2_f16[2];
  typedef i13 vec3_i13[3];

endpackage
