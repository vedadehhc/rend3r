`default_nettype none
`timescale 1ns / 1ps

import proctypes::*;

module fetch_tb;
    logic clk;
    logic rst;

    
    // 100 MHz clock
    always begin
        #5;
        clk = !clk;
    end

    FetchAction action;
    logic valid_out;
    InstructionAddr pc_out;
    Instruction inst_out;

    instruction_bank fetch (
        .clk(clk),
        .rst(rst),
        .action(action),
        .instruction_valid(valid_out),
        .pc_out(pc_out),
        .inst(inst_out)
    );

    initial begin
        $dumpfile("fetch.vcd");
        $dumpvars(0, fetch_tb);
        $display("Starting Sim");

        clk = 1'b0;
        rst = 1'b0;
        action = fetchStall;
        #10;
        #10;
        rst = 1'b1;
        #10;
        rst = 1'b0;
        #10;
        action = fetchDequeue;
        $display("");
        $display("Valid out: \t%32b", valid_out);
        $display("pc_out: \t%32b", pc_out);
        $display("inst_out \t%16b", inst_out);
        #10;
        action = fetchDequeue;
        $display("");
        $display("Valid out: \t%32b", valid_out);
        $display("pc_out: \t%32b", pc_out);
        $display("inst_out \t%16b", inst_out);
        #10;
        action = fetchDequeue;
        $display("");
        $display("Valid out: \t%32b", valid_out);
        $display("pc_out: \t%32b", pc_out);
        $display("inst_out \t%16b", inst_out);
        #10;
        action = fetchDequeue;
        $display("");
        $display("Valid out: \t%32b", valid_out);
        $display("pc_out: \t%32b", pc_out);
        $display("inst_out \t%16b", inst_out);
        #10;
        action = fetchDequeue;
        $display("");
        $display("Valid out: \t%32b", valid_out);
        $display("pc_out: \t%32b", pc_out);
        $display("inst_out \t%16b", inst_out);
        #10;
        action = fetchDequeue;
        $display("");
        $display("Valid out: \t%32b", valid_out);
        $display("pc_out: \t%32b", pc_out);
        $display("inst_out \t%16b", inst_out);
        #10;
        action = fetchDequeue;
        $display("");
        $display("Valid out: \t%32b", valid_out);
        $display("pc_out: \t%32b", pc_out);
        $display("inst_out \t%16b", inst_out);
        #10;
        action = fetchDequeue;
        $display("");
        $display("Valid out: \t%32b", valid_out);
        $display("pc_out: \t%32b", pc_out);
        $display("inst_out \t%16b", inst_out);
        #10;
        action = fetchDequeue;
        $display("");
        $display("Valid out: \t%32b", valid_out);
        $display("pc_out: \t%32b", pc_out);
        $display("inst_out \t%16b", inst_out);
        #10;
        action = fetchDequeue;
        $display("");
        $display("Valid out: \t%32b", valid_out);
        $display("pc_out: \t%32b", pc_out);
        $display("inst_out \t%16b", inst_out);
        #10;
        action = fetchDequeue;
        $display("");
        $display("Valid out: \t%32b", valid_out);
        $display("pc_out: \t%32b", pc_out);
        $display("inst_out \t%16b", inst_out);
        #10;
        action = fetchDequeue;
        $display("");
        $display("Valid out: \t%32b", valid_out);
        $display("pc_out: \t%32b", pc_out);
        $display("inst_out \t%16b", inst_out);
        #10;
        action = fetchDequeue;
        $display("");
        $display("Valid out: \t%32b", valid_out);
        $display("pc_out: \t%32b", pc_out);
        $display("inst_out \t%16b", inst_out);
        #10;
        action = fetchDequeue;
        $display("");
        $display("Valid out: \t%32b", valid_out);
        $display("pc_out: \t%32b", pc_out);
        $display("inst_out \t%16b", inst_out);
        #10;
        action = fetchDequeue;
        $display("");
        $display("Valid out: \t%32b", valid_out);
        $display("pc_out: \t%32b", pc_out);
        $display("inst_out \t%16b", inst_out);
        #10;
        action = fetchDequeue;
        $display("");
        $display("Valid out: \t%32b", valid_out);
        $display("pc_out: \t%32b", pc_out);
        $display("inst_out \t%16b", inst_out);
        #10;
        action = fetchDequeue;
        $display("");
        $display("Valid out: \t%32b", valid_out);
        $display("pc_out: \t%32b", pc_out);
        $display("inst_out \t%16b", inst_out);
        #10;
        action = fetchDequeue;
        $display("");
        $display("Valid out: \t%32b", valid_out);
        $display("pc_out: \t%32b", pc_out);
        $display("inst_out \t%16b", inst_out);

        #50;
        $display("\n\n");
        rst = 1'b0;
        action = fetchStall;
        #10;
        #10;
        rst = 1'b1;
        #10;
        rst = 1'b0;
        #30;
        action = fetchDequeue;
        $display("");
        $display("Valid out: \t%32b", valid_out);
        $display("pc_out: \t%32b", pc_out);
        $display("inst_out \t%16b", inst_out);
        #10;
        action = fetchStall;
        $display("");
        $display("Valid out: \t%32b", valid_out);
        $display("pc_out: \t%32b", pc_out);
        $display("inst_out \t%16b", inst_out);
        #10;
        action = fetchStall;
        $display("");
        $display("Valid out: \t%32b", valid_out);
        $display("pc_out: \t%32b", pc_out);
        $display("inst_out \t%16b", inst_out);
        #10;
        action = fetchStall;
        $display("");
        $display("Valid out: \t%32b", valid_out);
        $display("pc_out: \t%32b", pc_out);
        $display("inst_out \t%16b", inst_out);
        #10;
        action = fetchStall;
        $display("");
        $display("Valid out: \t%32b", valid_out);
        $display("pc_out: \t%32b", pc_out);
        $display("inst_out \t%16b", inst_out);
        #10;
        action = fetchDequeue;
        $display("");
        $display("Valid out: \t%32b", valid_out);
        $display("pc_out: \t%32b", pc_out);
        $display("inst_out \t%16b", inst_out);
        #10;
        action = fetchDequeue;
        $display("");
        $display("Valid out: \t%32b", valid_out);
        $display("pc_out: \t%32b", pc_out);
        $display("inst_out \t%16b", inst_out);
        #10;
        action = fetchDequeue;
        $display("");
        $display("Valid out: \t%32b", valid_out);
        $display("pc_out: \t%32b", pc_out);
        $display("inst_out \t%16b", inst_out);
        #10;
        action = fetchDequeue;
        $display("");
        $display("Valid out: \t%32b", valid_out);
        $display("pc_out: \t%32b", pc_out);
        $display("inst_out \t%16b", inst_out);
        #10;
        action = fetchDequeue;
        $display("");
        $display("Valid out: \t%32b", valid_out);
        $display("pc_out: \t%32b", pc_out);
        $display("inst_out \t%16b", inst_out);
        #10;
        action = fetchDequeue;
        $display("");
        $display("Valid out: \t%32b", valid_out);
        $display("pc_out: \t%32b", pc_out);
        $display("inst_out \t%16b", inst_out);
        #10;
        action = fetchDequeue;
        $display("");
        $display("Valid out: \t%32b", valid_out);
        $display("pc_out: \t%32b", pc_out);
        $display("inst_out \t%16b", inst_out);
        #10;
        action = fetchDequeue;
        $display("");
        $display("Valid out: \t%32b", valid_out);
        $display("pc_out: \t%32b", pc_out);
        $display("inst_out \t%16b", inst_out);
        #10;
        action = fetchDequeue;
        $display("");
        $display("Valid out: \t%32b", valid_out);
        $display("pc_out: \t%32b", pc_out);
        $display("inst_out \t%16b", inst_out);
        #10;
        action = fetchDequeue;
        $display("");
        $display("Valid out: \t%32b", valid_out);
        $display("pc_out: \t%32b", pc_out);
        $display("inst_out \t%16b", inst_out);
        #10;
        action = fetchDequeue;
        $display("");
        $display("Valid out: \t%32b", valid_out);
        $display("pc_out: \t%32b", pc_out);
        $display("inst_out \t%16b", inst_out);
        #10;
        action = fetchDequeue;
        $display("");
        $display("Valid out: \t%32b", valid_out);
        $display("pc_out: \t%32b", pc_out);
        $display("inst_out \t%16b", inst_out);
        #10;
        action = fetchDequeue;
        $display("");
        $display("Valid out: \t%32b", valid_out);
        $display("pc_out: \t%32b", pc_out);
        $display("inst_out \t%16b", inst_out);

        $display("\nFinishing Sim");
        $finish;
    end
endmodule